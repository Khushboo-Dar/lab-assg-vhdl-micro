version https://git-lfs.github.com/spec/v1
oid sha256:a489088c8ec93eaeed93d9f9e638be5ef5416d622551dbcb08f0f03af6c0dcac
size 925
