version https://git-lfs.github.com/spec/v1
oid sha256:4feb198e4acadb9790055d1a53f9e6de72f74f694e02ae34f47c40c681148cef
size 296
