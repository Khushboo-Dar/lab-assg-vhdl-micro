version https://git-lfs.github.com/spec/v1
oid sha256:afe5c239a63bfc5ac8f99599f48ef6f4899b0c3b07b88a1e02d1d5ac1d1b26b5
size 949
